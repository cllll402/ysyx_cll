module keycode_to_ascii(
    input [7:0] x,    
    output reg [7:0] y  
);
    always @(*) begin
        case (x)
            8'b00011100: y = 8'b01000001; // A 0x1C -> 0x41
            8'b00110010: y = 8'b01000010; // B 0x32 -> 0x42
            8'b00100001: y = 8'b01000011; // C 0x21 -> 0x43
            8'b00100011: y = 8'b01000100; // D 0x23 -> 0x44
            8'b00100100: y = 8'b01000101; // E 0x24 -> 0x45
            8'b00101011: y = 8'b01000110; // F 0x2B -> 0x46
            8'b00110100: y = 8'b01000111; // G 0x34 -> 0x47
            8'b00110011: y = 8'b01001000; // H 0x33 -> 0x48
            8'b01000011: y = 8'b01001001; // I 0x43 -> 0x49
            8'b00111011: y = 8'b01001010; // J 0x3B -> 0x4A
            8'b01000010: y = 8'b01001011; // K 0x42 -> 0x4B
            8'b01001011: y = 8'b01001100; // L 0x4B -> 0x4C
            8'b00111010: y = 8'b01001101; // M 0x3A -> 0x4D
            8'b00110001: y = 8'b01001110; // N 0x31 -> 0x4E
            8'b01000100: y = 8'b01001111; // O 0x44 -> 0x4F
            8'b01001101: y = 8'b01010000; // P 0x4D -> 0x50
            8'b00010101: y = 8'b01010001; // Q 0x15 -> 0x51
            8'b00101101: y = 8'b01010010; // R 0x2D -> 0x52
            8'b00011011: y = 8'b01010011; // S 0x1B -> 0x53
            8'b00101100: y = 8'b01010100; // T 0x2C -> 0x54
            8'b00111100: y = 8'b01010101; // U 0x3C -> 0x55
            8'b00101010: y = 8'b01010110; // V 0x2A -> 0x56
            8'b00011101: y = 8'b01010111; // W 0x1D -> 0x57
            8'b00100010: y = 8'b01011000; // X 0x22 -> 0x58
            8'b00110101: y = 8'b01011001; // Y 0x35 -> 0x59
            8'b00011010: y = 8'b01011010; // Z 0x1A -> 0x5A
            8'b01000101: y = 8'b00110000; // 0 0x45 -> 0x30
            8'b00010110: y = 8'b00110001; // 1 0x16 -> 0x31
            8'b00011110: y = 8'b00110010; // 2 0x1E -> 0x32
            8'b00100110: y = 8'b00110011; // 3 0x26 -> 0x33
            8'b00100101: y = 8'b00110100; // 4 0x25 -> 0x34
            8'b00101110: y = 8'b00110101; // 5 0x2E -> 0x35
            8'b00110110: y = 8'b00110110; // 6 0x36 -> 0x36
            8'b00111101: y = 8'b00110111; // 7 0x3D -> 0x37
            8'b00111110: y = 8'b00111000; // 8 0x3E -> 0x38
            8'b01000110: y = 8'b00111001; // 9 0x46 -> 0x39
            default: y = 8'b00000000;      
        endcase
    end
endmodule

