module bcd7hex(
	input [3:0] x,
	output reg [7:0] y
);
	
	always @ (*) begin 
		case (x)
			4'b0000 : y = 8'b00000010;  // 数码管显示 "0"
			4'b0001 : y = 8'b10011110;  // 数码管显示 "1"
			4'b0010 : y = 8'b00100100;  // 数码管显示 "2"
			4'b0011 : y = 8'b00001100;  // 数码管显示 "3"
			4'b0100 : y = 8'b10011000;  // 数码管显示 "4"
			4'b0101 : y = 8'b01001000;  // 数码管显示 "5"
			4'b0110 : y = 8'b01000000;  // 数码管显示 "6"
			4'b0111 : y = 8'b00011110;  // 数码管显示 "7"
			4'b1000 : y = 8'b00000000;  // 数码管显示 "8"
			4'b1001 : y = 8'b00001000;  // 数码管显示 "9"
			4'b1010 : y = 8'b00010000;  // 数码管显示 "A"
			4'b1011 : y = 8'b11000000;  // 数码管显示 "b"
			4'b1100 : y = 8'b01100010;  // 数码管显示 "C"
			4'b1101 : y = 8'b10000100;  // 数码管显示 "d"
			4'b1110 : y = 8'b01100000;  // 数码管显示 "E"
			4'b1111 : y = 8'b01110000;  // 数码管显示 "F"
			default : y = 8'b11111111;  // 默认全灭
		endcase
	end 
endmodule
	
	
